`timescale 1ns/1ns

//1- Module y Puertos 1/0
module ALUC (
		
		//Entradas
		input [2:0]OpA,
		input [5:0]Itr,
		
		//Salidas
		output reg [2:0]IA
);

//2- Delcaracion de señales --> NA(No aplica)

//3- Cuerpo del modulo

//Bloque Always
always @*

begin //Inicio_A	

	case (OpA)
		
		3'b000:
			
			case

				begin
				
			
				3'b000:



default:
	

endmodule