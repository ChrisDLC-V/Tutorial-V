module top_level (
    input [31:0] A,
    output reg R
);

endmodule //
